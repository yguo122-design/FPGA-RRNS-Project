`timescale 1ns / 1ps

module top_full_check(
    input wire clk,               // ��Ȼ���β�����Ҫ������߼���������ʱ�Ӷ˿�
    input wire [3:0] btn,         // BTN0 - BTN3
    
    // ��ɫ LED (LD4 - LD7)
    output wire [3:0] led,      
    
    // RGB LED LD0
    output wire led0_r, output wire led0_g, output wire led0_b,
    // RGB LED LD1
    output wire led1_r, output wire led1_g, output wire led1_b,
    // RGB LED LD2
    output wire led2_r, output wire led2_g, output wire led2_b,
    // RGB LED LD3
    output wire led3_r, output wire led3_g, output wire led3_b
    );

    // ------------------------------------------
    // 1. ��ɫ LED ���ԣ�ȫ������
    // ------------------------------------------
    assign led = 4'b1111;

    // ------------------------------------------
    // 2. RGB LED ��������
    // �߼���ÿ������һ��"Ĭ����ɫ"������Ӧ�İ�ť����ʱ���л���"������ɫ"
    // ------------------------------------------
    
    // --- LD0 ���� (��Ӧ BTN0) ---
    // Ĭ�ϣ���ɫ (R=1, G=0, B=0)
    // ���� BTN0����Ϊ ��ɫ (R=1, G=1, B=0) -> ֻ�� G ͨ���ܰ�ť����
    assign led0_r = 1'b1;
    assign led0_g = btn[0];       // ����(1)��ƣ��ɿ�(0)���
    assign led0_b = 1'b0;

    // --- LD1 ���� (��Ӧ BTN1) ---
    // Ĭ�ϣ���ɫ (R=0, G=1, B=0)
    // ���� BTN1����Ϊ ��ɫ (R=0, G=1, B=1) -> ֻ�� B ͨ���ܰ�ť����
    assign led1_r = 1'b0;
    assign led1_g = 1'b1;
    assign led1_b = btn[1];       // ����(1)���࣬�ɿ�(0)����

    // --- LD2 ���� (��Ӧ BTN2) ---
    // Ĭ�ϣ���ɫ (R=0, G=0, B=1)
    // ���� BTN2����Ϊ ��ɫ/Ʒ�� (R=1, G=0, B=1) -> ֻ�� R ͨ���ܰ�ť����
    assign led2_r = btn[2];       // ����(1)���ϣ��ɿ�(0)����
    assign led2_g = 1'b0;
    assign led2_b = 1'b1;

    // --- LD3 ���� (��Ӧ BTN3) ---
    // Ĭ�ϣ���ɫ (R=1, G=1, B=1)
    // ���� BTN3����Ϊ Ϩ�� (R=0, G=0, B=0) -> ����ͨ���ܰ�ť�������
    assign led3_r = ~btn[3];      // ����(1)��0(��)���ɿ�(0)��1(��)
    assign led3_g = ~btn[3];
    assign led3_b = ~btn[3];

endmodule